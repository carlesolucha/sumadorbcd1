library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--En realidad es un sumador de 4 bits normal y corriente
entity sumador4bits is 
	port(
	a : in std_logic_vector(3 downto 0);
	b : in std_logic_vector(3 downto 0);
	s : out std_logic_vector(3 downto 0);
	c_out : out std_logic);
end sumador4bits;

architecture structure of sumador4bits is
	signal c : std_logic_vector(4 downto 0);
	component sumador1
		port(
		a_i : in std_logic;
		b_i : in std_logic;
		c_i : in std_logic;
		s_i : out std_logic;
		c_i1 : out std_logic);
	end component;
begin
	c(0)<='0';
	c_out <= c(4);
	
	genSum : for i in 0 to 3 generate
	i_sumador4 : sumador1
		port map(
		a_i=>a(i),
		b_i=>b(i),
		s_i=>s(i),
		c_i=>c(i),
		c_i1=>c(i+1));
	end generate genSum;
end structure;